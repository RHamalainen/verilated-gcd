module tb_gcd;
endmodule
