module gcd (
    input clk,
    input rst,
    input in1,
    input in2,
    output out);

endmodule
